module equal_op(input a,input b,output result);
assign result=(a==b);
endmodule
