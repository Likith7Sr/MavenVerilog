module Left_Shift (  input [3:0] data,  output [7:0] result);
assign result = data << 2;
endmodule
